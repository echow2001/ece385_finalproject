////memory contents: to be filled in later. hard code to test data for cp1. 
//module memory_contents(input addr[10:0])
//    
//endmodule